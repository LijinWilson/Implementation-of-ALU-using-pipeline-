// --------- Pipeline modelling of an ALU ---------
// Here we are using non overlapping two phase clock


module pipeline_ALU(Zout, rs1, rs2, rd, func, addr,  clk1, clk2);
input [3:0] rs1, rs2, rd, func;
input [7:0] addr;
input clk1, clk2;

output [15:0] Zout;

// designing of intermediate storage elements
reg [15:0] L12_A, L12_B, L23_Z, L34_Z;
reg [3:0] L12_rd, L12_func, L23_rd;
reg [7:0] L12_addr, L23_addr, L34_addr;

// designing of register bank
reg [15:0] regBank [0:15];

// designing the memory element
reg [15:0] mem [0:255];

assign Zout = L34_Z;

// ------------- stage - 1 -------------
/*
 - In stage - 1 modelling we are inputting value of A and B
 - Forwarding the values of rd, func, addr;

*/

always @ (posedge clk1)
    begin
        L12_A <= #2 regBank[rs1];
        L12_B <= #2 regBank[rs2];
        L12_rd <= #2 rd;
        L12_func <= #2 func;
        L12_addr <= #2 addr;
    end

// ------------- stage - 2 -------------
    
always @ (negedge clk2)
    begin
        case(func)
            0: L23_Z <= #2  L12_A + L12_B; // addition
            1: L23_Z <= #2  L12_A - L12_B;
            2: L23_Z <= #2  L12_A * L12_B;
            3: L23_Z <= #2  L12_A;
            4: L23_Z <= #2  L12_B;
            5: L23_Z <= #2  L12_A & L12_B;
            6: L23_Z <= #2  L12_A | L12_B;
            7: L23_Z <= #2  L12_A ^ L12_B;
            8: L23_Z <= #2  ~L12_A;
            9: L23_Z <= #2  ~L12_B;
           10: L23_Z <= #2  L12_A >> 1;
           11: L23_Z <= #2  L12_A << 1;
           
           default: L23_Z <= #2 16'bxxxx;
        endcase
        
        L23_rd <= #2 L12_rd; 
        L23_addr <= #2 L12_addr;
        
    end
    
// ------------- stage - 3 -------------

always @ (posedge clk1)
    begin
        regBank[L23_rd] <= #2 L23_Z;
        L34_Z <= #2 L23_Z;
        L34_addr <= #2 L23_addr;
    end
    
// ------------- stage - 4 -------------
always @ (negedge clk2)
    begin
        mem[L34_addr] <= #2 L34_Z;
    end

endmodule

